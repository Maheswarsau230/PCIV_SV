module top;
initial begin
  $display("this is PCIE_SV");
end
endmodule
